
entity PIXELCODER is

end PIXELCODER;

architecture RTL of PIXELCODER is
begin

coder: process ()
begin

  case coderState is
  
    
  end case;
  
end process;

end RTL;